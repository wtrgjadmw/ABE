`define ALU_INST_BITS 42
`define MEM_SIZE 15
`define ADDR_BITS 4
`define CAL_MUX_BIT 2

`define INDEX_READA 0
`define INDEX_READB 7
`define INDEX_READC 14
`define INDEX_READD 20
`define INDEX_ISSUB 26
`define INDEX_MMVAL 27
`define INDEX_MASVAL 28
`define INDEX_WRITEA 29
`define INDEX_WRITEB 36
